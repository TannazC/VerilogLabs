module lab2part1 (SW, LEDR, HEX1, HEX0);
    //Initialize wires, LEDs, HEX (7seg)
    input [7:0] SW;
    output [7:0] LEDR;
    output [6:0] HEX1, HEX0;

    //wire [3:0] = s, c; not used here 
    assign LEDR[3:0] = SW[3:0];
    assign LEDR[7:4] = SW[7:4];

    //HEX0 7seg boolean eqns 
    assign HEX0[0] = (~SW[3]&~SW[2]&~SW[1]&SW[0])|(~SW[3]&SW[2]&~SW[1]&~SW[0]);
    assign HEX0[1] = (SW[2]&~SW[1]&SW[0])|(SW[2]&SW[1]&~SW[0]);
    assign HEX0[2] = (~SW[3]&~SW[2]&SW[1]&~SW[0]);
    assign HEX0[3] = (~SW[2]&~SW[1]&SW[0])|(SW[2]&~SW[1]&~SW[0])|(SW[2]&SW[1]&SW[0]);
    assign HEX0[4] = (SW[0])|(SW[2]&~SW[1]);
    assign HEX0[5] = (SW[1]&SW[0])|(~SW[2]&SW[1]&~SW[0])|(~SW[3]&~SW[2]&SW[0]);
    assign HEX0[6] = (~SW[3]&~SW[2]&~SW[1])|(SW[2]&SW[1]&SW[0]);

    //HEX1 7seg boolean eqns
    assign HEX1[0] = (~SW[7]&~SW[6]&~SW[5]&SW[4])|(~SW[7]&SW[6]&~SW[5]&~SW[4]);
    assign HEX1[1] = (SW[6]&~SW[5]&SW[4])|(SW[6]&SW[5]&~SW[4]);
    assign HEX1[2] = (~SW[7]&~SW[6]&SW[5]&~SW[4]);
    assign HEX1[3] = (~SW[6]&~SW[5]&SW[4])|(SW[6]&~SW[5]&~SW[4])|(SW[6]&SW[5]&SW[4]);
    assign HEX1[4] = (SW[4])|(SW[6]&~SW[5]);
    assign HEX1[5] = (SW[5]&SW[4])|(~SW[6]&SW[5]&~SW[4])|(~SW[7]&~SW[6]&SW[4]);
    assign HEX1[6] = (~SW[7]&~SW[6]&~SW[5])|(SW[6]&SW[5]&SW[4]);
endmodule